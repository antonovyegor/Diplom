library ieee;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;


entity test is 
end entity;

architecture SYN of test is 


begin


end SYN;