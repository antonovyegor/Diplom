CONV_INT_TO_FLOAT_inst : CONV_INT_TO_FLOAT PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
