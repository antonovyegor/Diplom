
module Debuger (
	source,
	probe);	

	output	[3:0]	source;
	input	[19:0]	probe;
endmodule
