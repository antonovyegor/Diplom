library ieee;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;



entity ROM12 is
	port (

			clock		: IN STD_LOGIC ;
			addr1		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q1		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr2		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q2		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr3		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q3		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr4		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q4		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr5		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q5		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr6		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q6		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr7		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q7		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr8		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q8		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr9		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q9		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr10		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q10		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr11		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q11		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			addr12		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			q12		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0)
			);
end entity;



architecture BEH of ROM12 is
subtype INT12 is  integer range 0 to 2047 ;
type MEM is array(0 to 1023) of INT12;
constant ROM : MEM :=(
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,1,1,1,
1,1,1,1,1,2,2,2,
2,2,2,2,3,3,3,3,
3,4,4,4,4,4,5,5,
5,5,6,6,6,6,7,7,
7,7,8,8,8,8,9,9,
9,10,10,10,11,11,11,12,
12,12,13,13,13,14,14,15,
15,15,16,16,16,17,17,18,
18,19,19,19,20,20,21,21,
22,22,23,23,24,24,25,25,
26,26,27,27,28,28,29,29,
30,30,31,31,32,32,33,34,
34,35,35,36,36,37,38,38,
39,39,40,41,41,42,43,43,
44,45,45,46,47,47,48,49,
49,50,51,51,52,53,53,54,
55,56,56,57,58,59,59,60,
61,62,62,63,64,65,66,66,
67,68,69,70,70,71,72,73,
74,75,75,76,77,78,79,80,
81,81,82,83,84,85,86,87,
88,89,89,90,91,92,93,94,
95,96,97,98,99,100,101,102,
103,104,105,106,107,108,109,110,
111,112,113,114,115,116,117,118,
119,120,121,122,123,125,126,127,
128,129,130,131,132,133,134,136,
137,138,139,140,141,142,144,145,
146,147,148,149,151,152,153,154,
155,157,158,159,160,161,163,164,
165,166,168,169,170,171,173,174,
175,176,178,179,180,182,183,184,
185,187,188,189,191,192,193,195,
196,197,199,200,201,203,204,206,
207,208,210,211,213,214,215,217,
218,220,221,222,224,225,227,228,
230,231,232,234,235,237,238,240,
241,243,244,246,247,249,250,252,
253,255,256,258,259,261,262,264,
265,267,269,270,272,273,275,276,
278,280,281,283,284,286,288,289,
291,292,294,296,297,299,301,302,
304,305,307,309,310,312,314,315,
317,319,321,322,324,326,327,329,
331,332,334,336,338,339,341,343,
345,346,348,350,352,353,355,357,
359,360,362,364,366,368,369,371,
373,375,377,378,380,382,384,386,
388,389,391,393,395,397,399,401,
402,404,406,408,410,412,414,416,
418,419,421,423,425,427,429,431,
433,435,437,439,441,443,445,446,
448,450,452,454,456,458,460,462,
464,466,468,470,472,474,476,478,
480,482,484,486,488,490,493,495,
497,499,501,503,505,507,509,511,
513,515,517,519,521,524,526,528,
530,532,534,536,538,540,543,545,
547,549,551,553,555,558,560,562,
564,566,568,571,573,575,577,579,
582,584,586,588,590,593,595,597,
599,601,604,606,608,610,613,615,
617,619,622,624,626,628,631,633,
635,637,640,642,644,647,649,651,
653,656,658,660,663,665,667,670,
672,674,677,679,681,684,686,688,
691,693,695,698,700,703,705,707,
710,712,714,717,719,722,724,726,
729,731,734,736,738,741,743,746,
748,751,753,755,758,760,763,765,
768,770,773,775,777,780,782,785,
787,790,792,795,797,800,802,805,
807,810,812,815,817,820,822,825,
827,830,832,835,837,840,842,845,
848,850,853,855,858,860,863,865,
868,871,873,876,878,881,883,886,
889,891,894,896,899,902,904,907,
909,912,915,917,920,923,925,928,
930,933,936,938,941,944,946,949,
952,954,957,960,962,965,968,970,
973,976,978,981,984,986,989,992,
994,997,1000,1002,1005,1008,1011,1013,
1016,1019,1021,1024,1027,1030,1032,1035,
1038,1041,1043,1046,1049,1051,1054,1057,
1060,1062,1065,1068,1071,1074,1076,1079,
1082,1085,1087,1090,1093,1096,1098,1101,
1104,1107,1110,1112,1115,1118,1121,1124,
1126,1129,1132,1135,1138,1140,1143,1146,
1149,1152,1155,1157,1160,1163,1166,1169,
1172,1174,1177,1180,1183,1186,1189,1192,
1194,1197,1200,1203,1206,1209,1212,1214,
1217,1220,1223,1226,1229,1232,1235,1237,
1240,1243,1246,1249,1252,1255,1258,1261,
1263,1266,1269,1272,1275,1278,1281,1284,
1287,1290,1293,1295,1298,1301,1304,1307,
1310,1313,1316,1319,1322,1325,1328,1331,
1334,1337,1340,1342,1345,1348,1351,1354,
1357,1360,1363,1366,1369,1372,1375,1378,
1381,1384,1387,1390,1393,1396,1399,1402,
1405,1408,1411,1414,1417,1420,1423,1426,
1429,1432,1435,1438,1441,1444,1447,1450,
1453,1456,1459,1462,1465,1468,1471,1474,
1477,1480,1483,1486,1489,1492,1495,1498,
1501,1504,1507,1510,1513,1516,1519,1522,
1525,1528,1531,1534,1537,1540,1543,1546,
1549,1553,1556,1559,1562,1565,1568,1571,
1574,1577,1580,1583,1586,1589,1592,1595,
1598,1601,1605,1608,1611,1614,1617,1620,
1623,1626,1629,1632,1635,1638,1641,1644,
1648,1651,1654,1657,1660,1663,1666,1669,
1672,1675,1678,1681,1685,1688,1691,1694,
1697,1700,1703,1706,1709,1712,1716,1719,
1722,1725,1728,1731,1734,1737,1740,1743,
1747,1750,1753,1756,1759,1762,1765,1768,
1771,1775,1778,1781,1784,1787,1790,1793,
1796,1799,1803,1806,1809,1812,1815,1818,
1821,1824,1828,1831,1834,1837,1840,1843,
1846,1849,1853,1856,1859,1862,1865,1868,
1871,1874,1878,1881,1884,1887,1890,1893,
1896,1900,1903,1906,1909,1912,1915,1918,
1921,1925,1928,1931,1934,1937,1940,1943,
1947,1950,1953,1956,1959,1962,1965,1968,
1972,1975,1978,1981,1984,1987,1990,1994,
1997,2000,2003,2006,2009,2012,2016,2019,
2022,2025,2028,2031,2034,2038,2041,2044--,


--2047,2050,2053,2056,2060,2063,2066,2069,
--2072,2075,2078,2082,2085,2088,2091,2094,
--2097,2100,2104,2107,2110,2113,2116,2119,
--2122,2126,2129,2132,2135,2138,2141,2144,
--2147,2151,2154,2157,2160,2163,2166,2169,
--2173,2176,2179,2182,2185,2188,2191,2194,
--2198,2201,2204,2207,2210,2213,2216,2220,
--2223,2226,2229,2232,2235,2238,2241,2245,
--2248,2251,2254,2257,2260,2263,2266,2270,
--2273,2276,2279,2282,2285,2288,2291,2295,
--2298,2301,2304,2307,2310,2313,2316,2319,
--2323,2326,2329,2332,2335,2338,2341,2344,
--2347,2351,2354,2357,2360,2363,2366,2369,
--2372,2375,2378,2382,2385,2388,2391,2394,
--2397,2400,2403,2406,2409,2413,2416,2419,
--2422,2425,2428,2431,2434,2437,2440,2443,
--2446,2450,2453,2456,2459,2462,2465,2468,
--2471,2474,2477,2480,2483,2486,2489,2493,
--2496,2499,2502,2505,2508,2511,2514,2517,
--2520,2523,2526,2529,2532,2535,2538,2541,
--2545,2548,2551,2554,2557,2560,2563,2566,
--2569,2572,2575,2578,2581,2584,2587,2590,
--2593,2596,2599,2602,2605,2608,2611,2614,
--2617,2620,2623,2626,2629,2632,2635,2638,
--2641,2644,2647,2650,2653,2656,2659,2662,
--2665,2668,2671,2674,2677,2680,2683,2686,
--2689,2692,2695,2698,2701,2704,2707,2710,
--2713,2716,2719,2722,2725,2728,2731,2734,
--2737,2740,2743,2746,2749,2752,2754,2757,
--2760,2763,2766,2769,2772,2775,2778,2781,
--2784,2787,2790,2793,2796,2799,2801,2804,
--2807,2810,2813,2816,2819,2822,2825,2828,
--2831,2833,2836,2839,2842,2845,2848,2851,
--2854,2857,2859,2862,2865,2868,2871,2874,
--2877,2880,2882,2885,2888,2891,2894,2897,
--2900,2902,2905,2908,2911,2914,2917,2920,
--2922,2925,2928,2931,2934,2937,2939,2942,
--2945,2948,2951,2954,2956,2959,2962,2965,
--2968,2970,2973,2976,2979,2982,2984,2987,
--2990,2993,2996,2998,3001,3004,3007,3009,
--3012,3015,3018,3020,3023,3026,3029,3032,
--3034,3037,3040,3043,3045,3048,3051,3053,
--3056,3059,3062,3064,3067,3070,3073,3075,
--3078,3081,3083,3086,3089,3092,3094,3097,
--3100,3102,3105,3108,3110,3113,3116,3118,
--3121,3124,3126,3129,3132,3134,3137,3140,
--3142,3145,3148,3150,3153,3156,3158,3161,
--3164,3166,3169,3171,3174,3177,3179,3182,
--3185,3187,3190,3192,3195,3198,3200,3203,
--3205,3208,3211,3213,3216,3218,3221,3223,
--3226,3229,3231,3234,3236,3239,3241,3244,
--3246,3249,3252,3254,3257,3259,3262,3264,
--3267,3269,3272,3274,3277,3279,3282,3284,
--3287,3289,3292,3294,3297,3299,3302,3304,
--3307,3309,3312,3314,3317,3319,3321,3324,
--3326,3329,3331,3334,3336,3339,3341,3343,
--3346,3348,3351,3353,3356,3358,3360,3363,
--3365,3368,3370,3372,3375,3377,3380,3382,
--3384,3387,3389,3391,3394,3396,3399,3401,
--3403,3406,3408,3410,3413,3415,3417,3420,
--3422,3424,3427,3429,3431,3434,3436,3438,
--3441,3443,3445,3447,3450,3452,3454,3457,
--3459,3461,3463,3466,3468,3470,3472,3475,
--3477,3479,3481,3484,3486,3488,3490,3493,
--3495,3497,3499,3501,3504,3506,3508,3510,
--3512,3515,3517,3519,3521,3523,3526,3528,
--3530,3532,3534,3536,3539,3541,3543,3545,
--3547,3549,3551,3554,3556,3558,3560,3562,
--3564,3566,3568,3570,3573,3575,3577,3579,
--3581,3583,3585,3587,3589,3591,3593,3595,
--3597,3599,3601,3604,3606,3608,3610,3612,
--3614,3616,3618,3620,3622,3624,3626,3628,
--3630,3632,3634,3636,3638,3640,3642,3644,
--3646,3648,3649,3651,3653,3655,3657,3659,
--3661,3663,3665,3667,3669,3671,3673,3675,
--3676,3678,3680,3682,3684,3686,3688,3690,
--3692,3693,3695,3697,3699,3701,3703,3705,
--3706,3708,3710,3712,3714,3716,3717,3719,
--3721,3723,3725,3726,3728,3730,3732,3734,
--3735,3737,3739,3741,3742,3744,3746,3748,
--3749,3751,3753,3755,3756,3758,3760,3762,
--3763,3765,3767,3768,3770,3772,3773,3775,
--3777,3779,3780,3782,3784,3785,3787,3789,
--3790,3792,3793,3795,3797,3798,3800,3802,
--3803,3805,3806,3808,3810,3811,3813,3814,
--3816,3818,3819,3821,3822,3824,3825,3827,
--3829,3830,3832,3833,3835,3836,3838,3839,
--3841,3842,3844,3845,3847,3848,3850,3851,
--3853,3854,3856,3857,3859,3860,3862,3863,
--3864,3866,3867,3869,3870,3872,3873,3874,
--3876,3877,3879,3880,3881,3883,3884,3886,
--3887,3888,3890,3891,3893,3894,3895,3897,
--3898,3899,3901,3902,3903,3905,3906,3907,
--3909,3910,3911,3912,3914,3915,3916,3918,
--3919,3920,3921,3923,3924,3925,3926,3928,
--3929,3930,3931,3933,3934,3935,3936,3937,
--3939,3940,3941,3942,3943,3945,3946,3947,
--3948,3949,3950,3952,3953,3954,3955,3956,
--3957,3958,3960,3961,3962,3963,3964,3965,
--3966,3967,3968,3969,3971,3972,3973,3974,
--3975,3976,3977,3978,3979,3980,3981,3982,
--3983,3984,3985,3986,3987,3988,3989,3990,
--3991,3992,3993,3994,3995,3996,3997,3998,
--3999,4000,4001,4002,4003,4004,4005,4005,
--4006,4007,4008,4009,4010,4011,4012,4013,
--4013,4014,4015,4016,4017,4018,4019,4019,
--4020,4021,4022,4023,4024,4024,4025,4026,
--4027,4028,4028,4029,4030,4031,4032,4032,
--4033,4034,4035,4035,4036,4037,4038,4038,
--4039,4040,4041,4041,4042,4043,4043,4044,
--4045,4045,4046,4047,4047,4048,4049,4049,
--4050,4051,4051,4052,4053,4053,4054,4055,
--4055,4056,4056,4057,4058,4058,4059,4059,
--4060,4060,4061,4062,4062,4063,4063,4064,
--4064,4065,4065,4066,4066,4067,4067,4068,
--4068,4069,4069,4070,4070,4071,4071,4072,
--4072,4073,4073,4074,4074,4075,4075,4075,
--4076,4076,4077,4077,4078,4078,4078,4079,
--4079,4079,4080,4080,4081,4081,4081,4082,
--4082,4082,4083,4083,4083,4084,4084,4084,
--4085,4085,4085,4086,4086,4086,4086,4087,
--4087,4087,4087,4088,4088,4088,4088,4089,
--4089,4089,4089,4090,4090,4090,4090,4090,
--4091,4091,4091,4091,4091,4092,4092,4092,
--4092,4092,4092,4092,4093,4093,4093,4093,
--4093,4093,4093,4093,4094,4094,4094,4094,
--4094,4094,4094,4094,4094,4094,4094,4094,
--4094,4094,4094,4094,4094,4094,4094,4094,
--4095,4094,4094,4094,4094,4094,4094,4094,
--4094,4094,4094,4094,4094,4094,4094,4094,
--4094,4094,4094,4094,4094,4093,4093,4093,
--4093,4093,4093,4093,4093,4092,4092,4092,
--4092,4092,4092,4092,4091,4091,4091,4091,
--4091,4090,4090,4090,4090,4090,4089,4089,
--4089,4089,4088,4088,4088,4088,4087,4087,
--4087,4087,4086,4086,4086,4086,4085,4085,
--4085,4084,4084,4084,4083,4083,4083,4082,
--4082,4082,4081,4081,4081,4080,4080,4079,
--4079,4079,4078,4078,4078,4077,4077,4076,
--4076,4075,4075,4075,4074,4074,4073,4073,
--4072,4072,4071,4071,4070,4070,4069,4069,
--4068,4068,4067,4067,4066,4066,4065,4065,
--4064,4064,4063,4063,4062,4062,4061,4060,
--4060,4059,4059,4058,4058,4057,4056,4056,
--4055,4055,4054,4053,4053,4052,4051,4051,
--4050,4049,4049,4048,4047,4047,4046,4045,
--4045,4044,4043,4043,4042,4041,4041,4040,
--4039,4038,4038,4037,4036,4035,4035,4034,
--4033,4032,4032,4031,4030,4029,4028,4028,
--4027,4026,4025,4024,4024,4023,4022,4021,
--4020,4019,4019,4018,4017,4016,4015,4014,
--4013,4013,4012,4011,4010,4009,4008,4007,
--4006,4005,4005,4004,4003,4002,4001,4000,
--3999,3998,3997,3996,3995,3994,3993,3992,
--3991,3990,3989,3988,3987,3986,3985,3984,
--3983,3982,3981,3980,3979,3978,3977,3976,
--3975,3974,3973,3972,3971,3969,3968,3967,
--3966,3965,3964,3963,3962,3961,3960,3958,
--3957,3956,3955,3954,3953,3952,3950,3949,
--3948,3947,3946,3945,3943,3942,3941,3940,
--3939,3937,3936,3935,3934,3933,3931,3930,
--3929,3928,3926,3925,3924,3923,3921,3920,
--3919,3918,3916,3915,3914,3912,3911,3910,
--3909,3907,3906,3905,3903,3902,3901,3899,
--3898,3897,3895,3894,3893,3891,3890,3888,
--3887,3886,3884,3883,3881,3880,3879,3877,
--3876,3874,3873,3872,3870,3869,3867,3866,
--3864,3863,3862,3860,3859,3857,3856,3854,
--3853,3851,3850,3848,3847,3845,3844,3842,
--3841,3839,3838,3836,3835,3833,3832,3830,
--3829,3827,3825,3824,3822,3821,3819,3818,
--3816,3814,3813,3811,3810,3808,3806,3805,
--3803,3802,3800,3798,3797,3795,3793,3792,
--3790,3789,3787,3785,3784,3782,3780,3779,
--3777,3775,3773,3772,3770,3768,3767,3765,
--3763,3762,3760,3758,3756,3755,3753,3751,
--3749,3748,3746,3744,3742,3741,3739,3737,
--3735,3734,3732,3730,3728,3726,3725,3723,
--3721,3719,3717,3716,3714,3712,3710,3708,
--3706,3705,3703,3701,3699,3697,3695,3693,
--3692,3690,3688,3686,3684,3682,3680,3678,
--3676,3675,3673,3671,3669,3667,3665,3663,
--3661,3659,3657,3655,3653,3651,3649,3648,
--3646,3644,3642,3640,3638,3636,3634,3632,
--3630,3628,3626,3624,3622,3620,3618,3616,
--3614,3612,3610,3608,3606,3604,3601,3599,
--3597,3595,3593,3591,3589,3587,3585,3583,
--3581,3579,3577,3575,3573,3570,3568,3566,
--3564,3562,3560,3558,3556,3554,3551,3549,
--3547,3545,3543,3541,3539,3536,3534,3532,
--3530,3528,3526,3523,3521,3519,3517,3515,
--3512,3510,3508,3506,3504,3501,3499,3497,
--3495,3493,3490,3488,3486,3484,3481,3479,
--3477,3475,3472,3470,3468,3466,3463,3461,
--3459,3457,3454,3452,3450,3447,3445,3443,
--3441,3438,3436,3434,3431,3429,3427,3424,
--3422,3420,3417,3415,3413,3410,3408,3406,
--3403,3401,3399,3396,3394,3391,3389,3387,
--3384,3382,3380,3377,3375,3372,3370,3368,
--3365,3363,3360,3358,3356,3353,3351,3348,
--3346,3343,3341,3339,3336,3334,3331,3329,
--3326,3324,3321,3319,3317,3314,3312,3309,
--3307,3304,3302,3299,3297,3294,3292,3289,
--3287,3284,3282,3279,3277,3274,3272,3269,
--3267,3264,3262,3259,3257,3254,3252,3249,
--3246,3244,3241,3239,3236,3234,3231,3229,
--3226,3223,3221,3218,3216,3213,3211,3208,
--3205,3203,3200,3198,3195,3192,3190,3187,
--3185,3182,3179,3177,3174,3171,3169,3166,
--3164,3161,3158,3156,3153,3150,3148,3145,
--3142,3140,3137,3134,3132,3129,3126,3124,
--3121,3118,3116,3113,3110,3108,3105,3102,
--3100,3097,3094,3092,3089,3086,3083,3081,
--3078,3075,3073,3070,3067,3064,3062,3059,
--3056,3053,3051,3048,3045,3043,3040,3037,
--3034,3032,3029,3026,3023,3020,3018,3015,
--3012,3009,3007,3004,3001,2998,2996,2993,
--2990,2987,2984,2982,2979,2976,2973,2970,
--2968,2965,2962,2959,2956,2954,2951,2948,
--2945,2942,2939,2937,2934,2931,2928,2925,
--2922,2920,2917,2914,2911,2908,2905,2902,
--2900,2897,2894,2891,2888,2885,2882,2880,
--2877,2874,2871,2868,2865,2862,2859,2857,
--2854,2851,2848,2845,2842,2839,2836,2833,
--2831,2828,2825,2822,2819,2816,2813,2810,
--2807,2804,2801,2799,2796,2793,2790,2787,
--2784,2781,2778,2775,2772,2769,2766,2763,
--2760,2757,2754,2752,2749,2746,2743,2740,
--2737,2734,2731,2728,2725,2722,2719,2716,
--2713,2710,2707,2704,2701,2698,2695,2692,
--2689,2686,2683,2680,2677,2674,2671,2668,
--2665,2662,2659,2656,2653,2650,2647,2644,
--2641,2638,2635,2632,2629,2626,2623,2620,
--2617,2614,2611,2608,2605,2602,2599,2596,
--2593,2590,2587,2584,2581,2578,2575,2572,
--2569,2566,2563,2560,2557,2554,2551,2548,
--2545,2541,2538,2535,2532,2529,2526,2523,
--2520,2517,2514,2511,2508,2505,2502,2499,
--2496,2493,2489,2486,2483,2480,2477,2474,
--2471,2468,2465,2462,2459,2456,2453,2450,
--2446,2443,2440,2437,2434,2431,2428,2425,
--2422,2419,2416,2413,2409,2406,2403,2400,
--2397,2394,2391,2388,2385,2382,2378,2375,
--2372,2369,2366,2363,2360,2357,2354,2351,
--2347,2344,2341,2338,2335,2332,2329,2326,
--2323,2319,2316,2313,2310,2307,2304,2301,
--2298,2295,2291,2288,2285,2282,2279,2276,
--2273,2270,2266,2263,2260,2257,2254,2251,
--2248,2245,2241,2238,2235,2232,2229,2226,
--2223,2220,2216,2213,2210,2207,2204,2201,
--2198,2194,2191,2188,2185,2182,2179,2176,
--2173,2169,2166,2163,2160,2157,2154,2151,
--2147,2144,2141,2138,2135,2132,2129,2126,
--2122,2119,2116,2113,2110,2107,2104,2100,
--2097,2094,2091,2088,2085,2082,2078,2075,
--2072,2069,2066,2063,2060,2056,2053,2050,
--2047,2044,2041,2038,2034,2031,2028,2025,
--2022,2019,2016,2012,2009,2006,2003,2000,
--1997,1994,1990,1987,1984,1981,1978,1975,
--1972,1968,1965,1962,1959,1956,1953,1950,
--1947,1943,1940,1937,1934,1931,1928,1925,
--1921,1918,1915,1912,1909,1906,1903,1900,
--1896,1893,1890,1887,1884,1881,1878,1874,
--1871,1868,1865,1862,1859,1856,1853,1849,
--1846,1843,1840,1837,1834,1831,1828,1824,
--1821,1818,1815,1812,1809,1806,1803,1799,
--1796,1793,1790,1787,1784,1781,1778,1775,
--1771,1768,1765,1762,1759,1756,1753,1750,
--1747,1743,1740,1737,1734,1731,1728,1725,
--1722,1719,1716,1712,1709,1706,1703,1700,
--1697,1694,1691,1688,1685,1681,1678,1675,
--1672,1669,1666,1663,1660,1657,1654,1651,
--1648,1644,1641,1638,1635,1632,1629,1626,
--1623,1620,1617,1614,1611,1608,1605,1601,
--1598,1595,1592,1589,1586,1583,1580,1577,
--1574,1571,1568,1565,1562,1559,1556,1553,
--1549,1546,1543,1540,1537,1534,1531,1528,
--1525,1522,1519,1516,1513,1510,1507,1504,
--1501,1498,1495,1492,1489,1486,1483,1480,
--1477,1474,1471,1468,1465,1462,1459,1456,
--1453,1450,1447,1444,1441,1438,1435,1432,
--1429,1426,1423,1420,1417,1414,1411,1408,
--1405,1402,1399,1396,1393,1390,1387,1384,
--1381,1378,1375,1372,1369,1366,1363,1360,
--1357,1354,1351,1348,1345,1342,1340,1337,
--1334,1331,1328,1325,1322,1319,1316,1313,
--1310,1307,1304,1301,1298,1295,1293,1290,
--1287,1284,1281,1278,1275,1272,1269,1266,
--1263,1261,1258,1255,1252,1249,1246,1243,
--1240,1237,1235,1232,1229,1226,1223,1220,
--1217,1214,1212,1209,1206,1203,1200,1197,
--1194,1192,1189,1186,1183,1180,1177,1174,
--1172,1169,1166,1163,1160,1157,1155,1152,
--1149,1146,1143,1140,1138,1135,1132,1129,
--1126,1124,1121,1118,1115,1112,1110,1107,
--1104,1101,1098,1096,1093,1090,1087,1085,
--1082,1079,1076,1074,1071,1068,1065,1062,
--1060,1057,1054,1051,1049,1046,1043,1041,
--1038,1035,1032,1030,1027,1024,1021,1019,
--1016,1013,1011,1008,1005,1002,1000,997,
--994,992,989,986,984,981,978,976,
--973,970,968,965,962,960,957,954,
--952,949,946,944,941,938,936,933,
--930,928,925,923,920,917,915,912,
--909,907,904,902,899,896,894,891,
--889,886,883,881,878,876,873,871,
--868,865,863,860,858,855,853,850,
--848,845,842,840,837,835,832,830,
--827,825,822,820,817,815,812,810,
--807,805,802,800,797,795,792,790,
--787,785,782,780,777,775,773,770,
--768,765,763,760,758,755,753,751,
--748,746,743,741,738,736,734,731,
--729,726,724,722,719,717,714,712,
--710,707,705,703,700,698,695,693,
--691,688,686,684,681,679,677,674,
--672,670,667,665,663,660,658,656,
--653,651,649,647,644,642,640,637,
--635,633,631,628,626,624,622,619,
--617,615,613,610,608,606,604,601,
--599,597,595,593,590,588,586,584,
--582,579,577,575,573,571,568,566,
--564,562,560,558,555,553,551,549,
--547,545,543,540,538,536,534,532,
--530,528,526,524,521,519,517,515,
--513,511,509,507,505,503,501,499,
--497,495,493,490,488,486,484,482,
--480,478,476,474,472,470,468,466,
--464,462,460,458,456,454,452,450,
--448,446,445,443,441,439,437,435,
--433,431,429,427,425,423,421,419,
--418,416,414,412,410,408,406,404,
--402,401,399,397,395,393,391,389,
--388,386,384,382,380,378,377,375,
--373,371,369,368,366,364,362,360,
--359,357,355,353,352,350,348,346,
--345,343,341,339,338,336,334,332,
--331,329,327,326,324,322,321,319,
--317,315,314,312,310,309,307,305,
--304,302,301,299,297,296,294,292,
--291,289,288,286,284,283,281,280,
--278,276,275,273,272,270,269,267,
--265,264,262,261,259,258,256,255,
--253,252,250,249,247,246,244,243,
--241,240,238,237,235,234,232,231,
--230,228,227,225,224,222,221,220,
--218,217,215,214,213,211,210,208,
--207,206,204,203,201,200,199,197,
--196,195,193,192,191,189,188,187,
--185,184,183,182,180,179,178,176,
--175,174,173,171,170,169,168,166,
--165,164,163,161,160,159,158,157,
--155,154,153,152,151,149,148,147,
--146,145,144,142,141,140,139,138,
--137,136,134,133,132,131,130,129,
--128,127,126,125,123,122,121,120,
--119,118,117,116,115,114,113,112,
--111,110,109,108,107,106,105,104,
--103,102,101,100,99,98,97,96,
--95,94,93,92,91,90,89,89,
--88,87,86,85,84,83,82,81,
--81,80,79,78,77,76,75,75,
--74,73,72,71,70,70,69,68,
--67,66,66,65,64,63,62,62,
--61,60,59,59,58,57,56,56,
--55,54,53,53,52,51,51,50,
--49,49,48,47,47,46,45,45,
--44,43,43,42,41,41,40,39,
--39,38,38,37,36,36,35,35,
--34,34,33,32,32,31,31,30,
--30,29,29,28,28,27,27,26,
--26,25,25,24,24,23,23,22,
--22,21,21,20,20,19,19,19,
--18,18,17,17,16,16,16,15,
--15,15,14,14,13,13,13,12,
--12,12,11,11,11,10,10,10,
--9,9,9,8,8,8,8,7,
--7,7,7,6,6,6,6,5,
--5,5,5,4,4,4,4,4,
--3,3,3,3,3,2,2,2,
--2,2,2,2,1,1,1,1,
--1,1,1,1,0,0,0,0,
--0,0,0,0,0,0,0,0,
--0,0,0,0,0,0,0,0
);
subtype addr is integer range 0 to 4095;



begin
		R1:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr1(11 downto 10) is 
					when "00" => addr:=addr1;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr1(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr1 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr1(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q1<=data;
				
				
				
			end if;
		end process;

		
		R2:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr2(11 downto 10) is 
					when "00" => addr:=addr2;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr2(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr2 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr2(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q2<=data;
				
				
				
			end if;
		end process;
		
		R3:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr3(11 downto 10) is 
					when "00" => addr:=addr3;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr3(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr3 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr3(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q3<=data;
				
				
				
			end if;
		end process;
		
		R4:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr4(11 downto 10) is 
					when "00" => addr:=addr4;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr4(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr4 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr4(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q4<=data;
				
				
				
			end if;
		end process;
		
		R5:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr5(11 downto 10) is 
					when "00" => addr:=addr5;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr5(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr5 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr5(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q5<=data;
				
				
				
			end if;
		end process;
		
		R6:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr6(11 downto 10) is 
					when "00" => addr:=addr6;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr6(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr6 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr6(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q6<=data;
				
				
				
			end if;
		end process;
		
		R7:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr7(11 downto 10) is 
					when "00" => addr:=addr7;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr7(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr7 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr7(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q7<=data;
				
				
				
			end if;
		end process;
		
		R8:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr8(11 downto 10) is 
					when "00" => addr:=addr8;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr8(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr8 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr8(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q8<=data;
				
				
				
			end if;
		end process;
		
		R9:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr9(11 downto 10) is 
					when "00" => addr:=addr9;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr9(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr9 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr9(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q9<=data;
				
				
				
			end if;
		end process;
		
		R10:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr10(11 downto 10) is 
					when "00" => addr:=addr10;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr10(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr10 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr10(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q10<=data;
				
				
				
			end if;
		end process;
		
		R11:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr11(11 downto 10) is 
					when "00" => addr:=addr11;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr11(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr11 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr11(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q11<=data;
				
				
				
			end if;
		end process;
		
		R12:process (clock)
		variable addr: std_LOGIC_VECTOR(11 downto 0 );
		variable data : std_LOGIC_VECTOR(11 downto 0 ) :=X"000" ;
		begin
			if (rising_edge(clock)) then
			
				case addr12(11 downto 10) is 
					when "00" => addr:=addr12;data:=conv_std_logic_vector (   ROM(conv_integer(addr))  , 12   );
					when "01" => addr:="00"& not(addr12(9 downto 0));data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "10" => addr:=addr12 xor X"800";data:=conv_std_logic_vector (  4095- ROM(conv_integer(addr))  , 12   );
					when "11" => addr:="00"& not(addr12(9 downto 0));
					when others => addr:=X"000";data:=conv_std_logic_vector (  ROM(conv_integer(addr))  , 12   ); 	
				end case;
				q12<=data;
				
				
				
			end if;
		end process;
		
		
		
	
end BEH;