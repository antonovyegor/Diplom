library ieee;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;



entity Block1 is 

port (
	C200: in std_LOGIC;
	C50 : in std_LOGIC;
	C10 : in std_LOGIC;
	ADDR : out std_LOGIC_VECTOR(11 dowNTO 0);
	DATA_SIN : in std_LOGIC_VECTOR(11 dowNTO 0);
	
	FREQ : in std_LOGIC_VECTOR(31 dowNTO 0) ;
	GATE : in std_LOGIC;
	MULT_OUT: in std_LOGIC_VECTOR (1 downto 0);
	BUSY : out std_LOGIC;
	
	ATTACK_TIME : in natural;
	DECAY_TIME : in natural;
	RELEASE_TIME : in natural;
		
	ATTACK_DELTA : in std_logic_vector(31 downto 0);
	DECAY_DELTA : in std_logic_vector(31 downto 0);
	RELEASE_DELTA : in std_logic_vector(31 downto 0);
		
	
	
	TO_ADD : out std_LOGIC_VECTOR(11 dowNTO 0)
);

end entity ;


architecture Syn of Block1 is 
	component Oscill 
		port (
			C: in std_logic;
			MULT_OUT : in std_LOGIC_VECTOR(1 downto 0);
			
			SIGNAL_OUT : out std_LOGIC_VECTOR (11 downto 0 );
			ADDRESS_OUT : out std_LOGIC_VECTOR (11 downto 0 );
			FROM_MEMORY : in  std_LOGIC_VECTOR (11 downto 0 );
			FREQ_REG : in std_logic_vector ( 31 downto 0 )

			);
	end component;
	component CONV_INT_TO_FLOAT
	port (
	clock : in std_logic;
	dataa : in std_LOGIC_VECTOR(12 downto 0);
	result: out std_LOGIC_VECTOR(31 downto 0)
	);
	end component;
	
	component MUL
	PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
	 end component;
	 
	 component CONV_FLOAT_TO_INT
	 port (
	clock : in std_logic;
	dataa : in std_LOGIC_VECTOR(31 downto 0);
	result: out std_LOGIC_VECTOR(12 downto 0)
	);
	end component;
	
	component ADSR
		port (
		C10 : in std_logic;
		C200 : in std_logic;
		R : in std_logic;
		GATE : in std_logic;
		BUSY : out std_logic;
		ATTACK_TIME : in natural;
		DECAY_TIME : in natural;
		RELEASE_TIME : in natural;
		
		ATTACK_DELTA : in std_logic_vector(31 downto 0);
		DECAY_DELTA : in std_logic_vector(31 downto 0);
		RELEASE_DELTA : in std_logic_vector(31 downto 0);
		
		FP : out std_logic_vector(31 downto 0)
		);
	end component;
	
	signal osc_out_int : std_LOGIC_VECTOR(12 dowNTO 0);
	signal osc_out_fp : std_LOGIC_VECTOR(31 dowNTO 0);
	signal mul_out_fp : std_LOGIC_VECTOR(31 dowNTO 0);
	signal mul_out_int : std_LOGIC_VECTOR(12 dowNTO 0);
	signal adsr_out_fp : std_LOGIC_VECTOR(31 dowNTO 0);

	
begin
	Oscill_inst : Oscill port map(C=>C50,MULT_OUT=>MULT_OUT,SIGNAL_OUT=>osc_out_int(11 downto 0),ADDRESS_OUT=>ADDR,FROM_MEMORY=>DATA_SIN,FREQ_REG=>FREQ);
	osc_out_int(12)<='0';
	
	
	
	CONV_INT_TO_FLOAT_inst : CONV_INT_TO_FLOAT PORT MAP (
		clock	 => C200,
		dataa	 => osc_out_int,
		result	 => osc_out_fp
	);
	
	
	MUL_inst : MUL port map (clock=>C200,dataa=>osc_out_fp,datab=>adsr_out_fp,result=>mul_out_fp);
	
	
	
	CONV_FLOAT_TO_INT_inst : CONV_FLOAT_TO_INT PORT MAP (
		clock	 => C200,
		dataa	 => mul_out_fp,
		result	 => mul_out_int
	);

	
	
	ADSR_inst: ADSR port map(FP=>adsr_out_fp,c200=>c200,C10=>c10,R=>'0',gatE=>GATE,busy=>BUSY,attACK_TIME=>ATTACK_TIME,decAY_TIME=>DECAY_TIME,relEASE_TIME=>RELEASE_TIME,attACK_DELTA=>ATTACK_DELTA,decAY_DELTA=>DECAY_DELTA,
	relEASE_DELTA=>relEASE_DELTA);
	
	TO_ADD<=mul_out_int(11 downto 0);
end Syn;