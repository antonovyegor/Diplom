CONV_FLOAT_TO_INT_inst : CONV_FLOAT_TO_INT PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
