-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
-- CREATED		"Thu Jun 13 16:40:25 2019"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 



ENTITY MAINDIAGRAM IS 
	PORT
	(
		C :  IN  STD_LOGIC;
		R :  IN  STD_LOGIC;
		RX :  IN  STD_LOGIC;
		BUT1 :  IN  STD_LOGIC;
		BUT2 :  IN  STD_LOGIC;
		BUTTONS :  IN  STD_LOGIC_VECTOR(0 TO 11);
		SIGNAL_OUT :  OUT  STD_LOGIC
	);
END MAINDIAGRAM;

ARCHITECTURE bdf_type OF MAINDIAGRAM IS 

COMPONENT block1
	PORT(C200 : IN STD_LOGIC;
		 C50 : IN STD_LOGIC;
		 C10 : IN STD_LOGIC;
		 GATE : IN STD_LOGIC;
		 ATTACK_DELTA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ATTACK_TIME : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
		 DATA_SIN : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 DECAY_DELTA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DECAY_TIME : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
		 FREQ : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MULT_OUT : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 RELEASE_DELTA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RELEASE_TIME : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
		 BUSY : OUT STD_LOGIC;
		 ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		 TO_ADD : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dac
	PORT(DAC_Clk : IN STD_LOGIC;
		 DACin : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
		 DACout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT add
	PORT(data0x : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
	);
END COMPONENT;

COMPONENT romserial
	PORT(clock400 : IN STD_LOGIC;
		 addr0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 addr1 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 data0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		 data1 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pll
	PORT(inclk0 : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 c1 : OUT STD_LOGIC;
		 c2 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT buttonproc
	PORT(C200 : IN STD_LOGIC;
		 BUSY1 : IN STD_LOGIC;
		 BUSY2 : IN STD_LOGIC;
		 BUTTON : IN STD_LOGIC_VECTOR(0 TO 11);
		 OCTAVE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 GATE1 : OUT STD_LOGIC;
		 GATE2 : OUT STD_LOGIC;
		 FREQ1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FREQ2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uartproc
	PORT(C : IN STD_LOGIC;
		 R : IN STD_LOGIC;
		 READY : IN STD_LOGIC;
		 BUT_1 : IN STD_LOGIC;
		 BUT_2 : IN STD_LOGIC;
		 DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ATTACK_DELTA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ATTACK_TIME : OUT STD_LOGIC_VECTOR(30 DOWNTO 0);
		 DECAY_DELTA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DECAY_TIME : OUT STD_LOGIC_VECTOR(30 DOWNTO 0);
		 MULT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 OCTAVE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 RELEASE_DELTA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RELEASE_TIME : OUT STD_LOGIC_VECTOR(30 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uartrx
	PORT(clk50 : IN STD_LOGIC;
		 R : IN STD_LOGIC;
		 RX : IN STD_LOGIC;
		 ready : OUT STD_LOGIC;
		 RXOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(30 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(30 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(30 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(12 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(7 DOWNTO 0);


BEGIN 



b2v_inst : block1
PORT MAP(C200 => SYNTHESIZED_WIRE_37,
		 C50 => C,
		 C10 => SYNTHESIZED_WIRE_38,
		 GATE => SYNTHESIZED_WIRE_2,
		 ATTACK_DELTA => SYNTHESIZED_WIRE_39,
		 ATTACK_TIME => SYNTHESIZED_WIRE_40,
		 DATA_SIN => SYNTHESIZED_WIRE_5,
		 DECAY_DELTA => SYNTHESIZED_WIRE_41,
		 DECAY_TIME => SYNTHESIZED_WIRE_42,
		 FREQ => SYNTHESIZED_WIRE_8,
		 MULT_OUT => SYNTHESIZED_WIRE_43,
		 RELEASE_DELTA => SYNTHESIZED_WIRE_44,
		 RELEASE_TIME => SYNTHESIZED_WIRE_45,
		 BUSY => SYNTHESIZED_WIRE_31,
		 ADDR => SYNTHESIZED_WIRE_28,
		 TO_ADD => SYNTHESIZED_WIRE_26);


b2v_inst1 : dac
PORT MAP(DAC_Clk => C,
		 DACin => SYNTHESIZED_WIRE_12,
		 DACout => SIGNAL_OUT);


b2v_inst11 : block1
PORT MAP(C200 => SYNTHESIZED_WIRE_37,
		 C50 => C,
		 C10 => SYNTHESIZED_WIRE_38,
		 GATE => SYNTHESIZED_WIRE_15,
		 ATTACK_DELTA => SYNTHESIZED_WIRE_39,
		 ATTACK_TIME => SYNTHESIZED_WIRE_40,
		 DATA_SIN => SYNTHESIZED_WIRE_18,
		 DECAY_DELTA => SYNTHESIZED_WIRE_41,
		 DECAY_TIME => SYNTHESIZED_WIRE_42,
		 FREQ => SYNTHESIZED_WIRE_21,
		 MULT_OUT => SYNTHESIZED_WIRE_43,
		 RELEASE_DELTA => SYNTHESIZED_WIRE_44,
		 RELEASE_TIME => SYNTHESIZED_WIRE_45,
		 BUSY => SYNTHESIZED_WIRE_32,
		 ADDR => SYNTHESIZED_WIRE_29,
		 TO_ADD => SYNTHESIZED_WIRE_25);


b2v_inst12 : add
PORT MAP(data0x => SYNTHESIZED_WIRE_25,
		 data1x => SYNTHESIZED_WIRE_26,
		 result => SYNTHESIZED_WIRE_12);


b2v_inst2 : romserial
PORT MAP(clock400 => SYNTHESIZED_WIRE_37,
		 addr0 => SYNTHESIZED_WIRE_28,
		 addr1 => SYNTHESIZED_WIRE_29,
		 data0 => SYNTHESIZED_WIRE_5,
		 data1 => SYNTHESIZED_WIRE_18);


b2v_inst3 : pll
PORT MAP(inclk0 => C,
		 c0 => SYNTHESIZED_WIRE_46,
		 c1 => SYNTHESIZED_WIRE_37,
		 c2 => SYNTHESIZED_WIRE_38);


b2v_inst7 : buttonproc
PORT MAP(C200 => SYNTHESIZED_WIRE_46,
		 BUSY1 => SYNTHESIZED_WIRE_31,
		 BUSY2 => SYNTHESIZED_WIRE_32,
		 BUTTON => BUTTONS,
		 OCTAVE => SYNTHESIZED_WIRE_33,
		 GATE1 => SYNTHESIZED_WIRE_2,
		 GATE2 => SYNTHESIZED_WIRE_15,
		 FREQ1 => SYNTHESIZED_WIRE_8,
		 FREQ2 => SYNTHESIZED_WIRE_21);


b2v_inst8 : uartproc
PORT MAP(C => SYNTHESIZED_WIRE_46,
		 R => R,
		 READY => SYNTHESIZED_WIRE_35,
		 BUT_1 => BUT1,
		 BUT_2 => BUT2,
		 DATA => SYNTHESIZED_WIRE_36,
		 ATTACK_DELTA => SYNTHESIZED_WIRE_39,
		 ATTACK_TIME => SYNTHESIZED_WIRE_40,
		 DECAY_DELTA => SYNTHESIZED_WIRE_41,
		 DECAY_TIME => SYNTHESIZED_WIRE_42,
		 MULT => SYNTHESIZED_WIRE_43,
		 OCTAVE => SYNTHESIZED_WIRE_33,
		 RELEASE_DELTA => SYNTHESIZED_WIRE_44,
		 RELEASE_TIME => SYNTHESIZED_WIRE_45);


b2v_inst9 : uartrx
PORT MAP(clk50 => C,
		 R => R,
		 RX => RX,
		 ready => SYNTHESIZED_WIRE_35,
		 RXOUT => SYNTHESIZED_WIRE_36);


END bdf_type;